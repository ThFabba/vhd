conectix             0�{win   Wi2k     0       0   Z   ���D�A4��3�B��/Tp�+                                                                                                                                                                                                                                                                                                                                                                                                                                             cxsparse��������                 ���u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        conectix             0�{win   Wi2k     0       0   Z   ���D�A4��3�B��/Tp�+                                                                                                                                                                                                                                                                                                                                                                                                                                             